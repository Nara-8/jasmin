(** This module is meant as the minimal dependency of extracted code. *)
Require compiler.
Require psem_defs.
Require arm_params.
Require x86_params.
Require riscv_params.
Require sem_params_of_arch_extra.
Require wint_to_int.
